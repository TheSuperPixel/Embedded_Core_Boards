//****************************************Copyright (c)***********************************//
//ԭ�Ӹ����߽�ѧƽ̨��www.yuanzige.com
//����֧�֣�http://www.openedv.com/forum.php
//�Ա����̣�https://zhengdianyuanzi.tmall.com
//��ע΢�Ź���ƽ̨΢�źţ�"����ԭ��"����ѻ�ȡZYNQ & FPGA & STM32 & LINUX���ϡ�
//��Ȩ���У�����ؾ���
//Copyright(C) ����ԭ�� 2023-2033
//All rights reserved                                  
//----------------------------------------------------------------------------------------
// File name:           key_led
// Created by:          ����ԭ��
// Created date:        2023��2��22��14:17:02
// Version:             V1.0
// Descriptions:        ��������LED��ʵ��
//
//----------------------------------------------------------------------------------------
//****************************************************************************************//
module key_led(
    //input
    input               sys_clk,
    input               sys_rst_n,
    input        [4:0]  key,
    //output        
    output  reg  [4:0]  led 
    );

ila_0 key_ila_0 (
	.clk(sys_clk), // input wire clk


	.probe0(key) // input wire [4:0] probe0
);
//����
parameter CNT_MAX = 25'd25000000;    

//reg define
reg  [24:0]  cnt;
reg  [1:0]   led_flag;

//*****************************************************
//**                    main code
//*****************************************************

//��������ʱ0.5s
always @(posedge sys_clk or negedge sys_rst_n) begin
    if(!sys_rst_n)
        cnt <= 25'd0;
    else if(cnt < (CNT_MAX - 25'd1))
        cnt <= cnt + 25'd1;
    else
        cnt <= 25'd0;
end

//LED״̬�л���־λ
//  0  1  2  3
//  00 01 10 11
always @(posedge sys_clk or negedge sys_rst_n) begin
    if(!sys_rst_n)
        led_flag <= 2'd0;
    else if(cnt == (CNT_MAX - 25'd1))   
        led_flag <= led_flag + 2'd1;
    else
        led_flag <= led_flag;
end    
    
//LED����(�����ĸ�KEY�����£���led_flag����LED���и�ֵ)
always @(posedge sys_clk or negedge sys_rst_n) begin
    if(!sys_rst_n)
        led <= 5'b0000;
    else begin
        case(key)
            5'b11111 : led <= 5'b0000;
            5'b11110 : begin 
                if(led_flag == 2'd0)
                    led <= 5'b00001;
                else
                    led <= 5'b00000; 
            end
            5'b11101 : begin 
                if(led_flag == 2'd0)
                    led <= 5'b00010;
                else
                    led <= 5'b00000; 
            end  
            5'b11011 : begin 
                if(led_flag == 2'd0)
                    led <= 5'b00100;
                else
                    led <= 5'b00000; 
            end        
            5'b10111 : begin
                if(led_flag == 2'd0)
                    led <= 5'b01000;
                else
                    led <= 5'b00000; 
            end
            5'b01111 : begin
                if(led_flag == 2'd0)
                    led <= 5'b10000;
                else
                    led <= 5'b00000; 
            end
            default : ;
        endcase    
    end
end      
    
endmodule
